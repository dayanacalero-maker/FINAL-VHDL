library verilog;
use verilog.vl_types.all;
entity TOP_ALU_vlg_vec_tst is
end TOP_ALU_vlg_vec_tst;
